----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Twsa Liu
-- 
-- Create Date:    14:35:22 07/28/2017 
-- Design Name: 
-- Module Name:    multiplex_4_to_1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: ��ѡһ��·ѡ����VHDLģ�ͼ�����ƽ̨
--
-- Dependencies:  
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity multiplex_4_to_1 is
    Port ( 
	        clk :in STD_LOGIC;
	        a : in  STD_LOGIC_VECTOR (3 downto 0);
           sel : in  STD_LOGIC_VECTOR (1 downto 0);
           z : out  STD_LOGIC);
end multiplex_4_to_1;

architecture eqn of multiplex_4_to_1 is

begin
   with sel select
	z <= a(0) when "00",
	     a(1) when "01",
        a(2) when "10",
	     a(3) when others;
	
end architecture eqn;

